`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/11/30 19:38:34
// Design Name: 
// Module Name: ALU_Control
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ALU_Control(
    input [3:0] ALUOp,//�����źţ�ALU�ֲ�����
    input [5:0] func,//R��ָ���function��
    
    output reg ALUSrcA, ALUSrcB,//���ALU����ѡ���ź�
    output reg [2:0] ALUCtr//ALU�������
    );
    
    //ALU�ֲ�����
    always @ (*) begin
        if (ALUOp[3] == 1) begin
            ALUSrcA = (func == 6'b000000) ? 1 : 0;
            ALUSrcB = 0;
            ALUCtr[2] = (func == 6'b000000) ? 1 : 0;
            ALUCtr[1] = (func == 6'b100100 || func == 6'b100101) ? 1 : 0;
            ALUCtr[0] = (func == 6'b100010 || func == 6'b100101) ? 1 : 0;
        end
        else begin
            ALUSrcA = 0;
            ALUSrcB = (ALUOp == 4'b0001) ? 0 : 1;
            ALUCtr[2] = (ALUOp == 4'b0101 || ALUOp == 4'b0110) ? 1 : 0;
            ALUCtr[1] = (ALUOp == 4'b0010 || ALUOp == 4'b0011 || ALUOp == 4'b0110) ? 1 : 0;
            ALUCtr[0] = (ALUOp == 4'b0011 || ALUOp == 4'b0101 || ALUOp == 4'b0001) ? 1 : 0;
        end
    end
    
endmodule
