`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/12/09 18:08:22
// Design Name: 
// Module Name: Transfer
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Transfer(
    input CLK,//��Ƶ���ʱ��
    input [15:0] In,//������Ҫ��ʾ������
    
    output reg [3:0] Out,//��Ҫ��ʾ��������ϵ����֣�1λ��
    output reg [3:0] Bit//�����ɨ���ź�
    );

//���ڱ�����Ҫ��ʾ���źŵ�ÿһλ����Ӧ����Ե������
integer i;
initial begin
    i = 0;
end

//ѡ����Ҫ��ʾ�����ݺ���Ҫ�����������
always @ (negedge CLK) begin
    case(i)
        0 : begin
            Out = In [15:12];
            Bit = 4'b1110;
        end
        1 : begin
            Out = In [11:8];
            Bit = 4'b1101;
        end
        2 : begin
            Out = In [7:4];
            Bit = 4'b1011;
        end
        3 : begin
            Out = In [3:0];
            Bit = 4'b0111;
        end
    endcase
    i = (i == 3) ? 0 : i + 1;
end

endmodule
